module costable (
	input wire [9:0] cnt,
	output wire [9:0] cv
);

assign cv = cos(cnt);

function [9:0] cos(input[9:0] inp);
	begin
		case(inp)
		10'd   0: cos = 10'd1023;
		10'd   1: cos = 10'd1022;
		10'd   2: cos = 10'd1022;
		10'd   3: cos = 10'd1022;
		10'd   4: cos = 10'd1022;
		10'd   5: cos = 10'd1022;
		10'd   6: cos = 10'd1022;
		10'd   7: cos = 10'd1022;
		10'd   8: cos = 10'd1022;
		10'd   9: cos = 10'd1022;
		10'd  10: cos = 10'd1022;
		10'd  11: cos = 10'd1021;
		10'd  12: cos = 10'd1021;
		10'd  13: cos = 10'd1021;
		10'd  14: cos = 10'd1021;
		10'd  15: cos = 10'd1020;
		10'd  16: cos = 10'd1020;
		10'd  17: cos = 10'd1020;
		10'd  18: cos = 10'd1019;
		10'd  19: cos = 10'd1019;
		10'd  20: cos = 10'd1019;
		10'd  21: cos = 10'd1018;
		10'd  22: cos = 10'd1018;
		10'd  23: cos = 10'd1017;
		10'd  24: cos = 10'd1017;
		10'd  25: cos = 10'd1016;
		10'd  26: cos = 10'd1016;
		10'd  27: cos = 10'd1015;
		10'd  28: cos = 10'd1015;
		10'd  29: cos = 10'd1014;
		10'd  30: cos = 10'd1014;
		10'd  31: cos = 10'd1013;
		10'd  32: cos = 10'd1013;
		10'd  33: cos = 10'd1012;
		10'd  34: cos = 10'd1011;
		10'd  35: cos = 10'd1011;
		10'd  36: cos = 10'd1010;
		10'd  37: cos = 10'd1009;
		10'd  38: cos = 10'd1009;
		10'd  39: cos = 10'd1008;
		10'd  40: cos = 10'd1007;
		10'd  41: cos = 10'd1006;
		10'd  42: cos = 10'd1006;
		10'd  43: cos = 10'd1005;
		10'd  44: cos = 10'd1004;
		10'd  45: cos = 10'd1003;
		10'd  46: cos = 10'd1002;
		10'd  47: cos = 10'd1001;
		10'd  48: cos = 10'd1000;
		10'd  49: cos = 10'd1000;
		10'd  50: cos = 10'd999;
		10'd  51: cos = 10'd998;
		10'd  52: cos = 10'd997;
		10'd  53: cos = 10'd996;
		10'd  54: cos = 10'd995;
		10'd  55: cos = 10'd994;
		10'd  56: cos = 10'd993;
		10'd  57: cos = 10'd992;
		10'd  58: cos = 10'd990;
		10'd  59: cos = 10'd989;
		10'd  60: cos = 10'd988;
		10'd  61: cos = 10'd987;
		10'd  62: cos = 10'd986;
		10'd  63: cos = 10'd985;
		10'd  64: cos = 10'd984;
		10'd  65: cos = 10'd982;
		10'd  66: cos = 10'd981;
		10'd  67: cos = 10'd980;
		10'd  68: cos = 10'd979;
		10'd  69: cos = 10'd977;
		10'd  70: cos = 10'd976;
		10'd  71: cos = 10'd975;
		10'd  72: cos = 10'd973;
		10'd  73: cos = 10'd972;
		10'd  74: cos = 10'd971;
		10'd  75: cos = 10'd969;
		10'd  76: cos = 10'd968;
		10'd  77: cos = 10'd966;
		10'd  78: cos = 10'd965;
		10'd  79: cos = 10'd964;
		10'd  80: cos = 10'd962;
		10'd  81: cos = 10'd961;
		10'd  82: cos = 10'd959;
		10'd  83: cos = 10'd958;
		10'd  84: cos = 10'd956;
		10'd  85: cos = 10'd954;
		10'd  86: cos = 10'd953;
		10'd  87: cos = 10'd951;
		10'd  88: cos = 10'd950;
		10'd  89: cos = 10'd948;
		10'd  90: cos = 10'd946;
		10'd  91: cos = 10'd945;
		10'd  92: cos = 10'd943;
		10'd  93: cos = 10'd941;
		10'd  94: cos = 10'd940;
		10'd  95: cos = 10'd938;
		10'd  96: cos = 10'd936;
		10'd  97: cos = 10'd935;
		10'd  98: cos = 10'd933;
		10'd  99: cos = 10'd931;
		10'd 100: cos = 10'd929;
		10'd 101: cos = 10'd927;
		10'd 102: cos = 10'd926;
		10'd 103: cos = 10'd924;
		10'd 104: cos = 10'd922;
		10'd 105: cos = 10'd920;
		10'd 106: cos = 10'd918;
		10'd 107: cos = 10'd916;
		10'd 108: cos = 10'd914;
		10'd 109: cos = 10'd912;
		10'd 110: cos = 10'd910;
		10'd 111: cos = 10'd908;
		10'd 112: cos = 10'd906;
		10'd 113: cos = 10'd904;
		10'd 114: cos = 10'd902;
		10'd 115: cos = 10'd900;
		10'd 116: cos = 10'd898;
		10'd 117: cos = 10'd896;
		10'd 118: cos = 10'd894;
		10'd 119: cos = 10'd892;
		10'd 120: cos = 10'd890;
		10'd 121: cos = 10'd888;
		10'd 122: cos = 10'd886;
		10'd 123: cos = 10'd884;
		10'd 124: cos = 10'd881;
		10'd 125: cos = 10'd879;
		10'd 126: cos = 10'd877;
		10'd 127: cos = 10'd875;
		10'd 128: cos = 10'd873;
		10'd 129: cos = 10'd870;
		10'd 130: cos = 10'd868;
		10'd 131: cos = 10'd866;
		10'd 132: cos = 10'd864;
		10'd 133: cos = 10'd861;
		10'd 134: cos = 10'd859;
		10'd 135: cos = 10'd857;
		10'd 136: cos = 10'd855;
		10'd 137: cos = 10'd852;
		10'd 138: cos = 10'd850;
		10'd 139: cos = 10'd847;
		10'd 140: cos = 10'd845;
		10'd 141: cos = 10'd843;
		10'd 142: cos = 10'd840;
		10'd 143: cos = 10'd838;
		10'd 144: cos = 10'd835;
		10'd 145: cos = 10'd833;
		10'd 146: cos = 10'd831;
		10'd 147: cos = 10'd828;
		10'd 148: cos = 10'd826;
		10'd 149: cos = 10'd823;
		10'd 150: cos = 10'd821;
		10'd 151: cos = 10'd818;
		10'd 152: cos = 10'd816;
		10'd 153: cos = 10'd813;
		10'd 154: cos = 10'd811;
		10'd 155: cos = 10'd808;
		10'd 156: cos = 10'd806;
		10'd 157: cos = 10'd803;
		10'd 158: cos = 10'd800;
		10'd 159: cos = 10'd798;
		10'd 160: cos = 10'd795;
		10'd 161: cos = 10'd793;
		10'd 162: cos = 10'd790;
		10'd 163: cos = 10'd787;
		10'd 164: cos = 10'd785;
		10'd 165: cos = 10'd782;
		10'd 166: cos = 10'd779;
		10'd 167: cos = 10'd777;
		10'd 168: cos = 10'd774;
		10'd 169: cos = 10'd771;
		10'd 170: cos = 10'd769;
		10'd 171: cos = 10'd766;
		10'd 172: cos = 10'd763;
		10'd 173: cos = 10'd760;
		10'd 174: cos = 10'd758;
		10'd 175: cos = 10'd755;
		10'd 176: cos = 10'd752;
		10'd 177: cos = 10'd749;
		10'd 178: cos = 10'd747;
		10'd 179: cos = 10'd744;
		10'd 180: cos = 10'd741;
		10'd 181: cos = 10'd738;
		10'd 182: cos = 10'd735;
		10'd 183: cos = 10'd733;
		10'd 184: cos = 10'd730;
		10'd 185: cos = 10'd727;
		10'd 186: cos = 10'd724;
		10'd 187: cos = 10'd721;
		10'd 188: cos = 10'd718;
		10'd 189: cos = 10'd715;
		10'd 190: cos = 10'd713;
		10'd 191: cos = 10'd710;
		10'd 192: cos = 10'd707;
		10'd 193: cos = 10'd704;
		10'd 194: cos = 10'd701;
		10'd 195: cos = 10'd698;
		10'd 196: cos = 10'd695;
		10'd 197: cos = 10'd692;
		10'd 198: cos = 10'd689;
		10'd 199: cos = 10'd686;
		10'd 200: cos = 10'd683;
		10'd 201: cos = 10'd680;
		10'd 202: cos = 10'd677;
		10'd 203: cos = 10'd674;
		10'd 204: cos = 10'd671;
		10'd 205: cos = 10'd668;
		10'd 206: cos = 10'd665;
		10'd 207: cos = 10'd662;
		10'd 208: cos = 10'd659;
		10'd 209: cos = 10'd656;
		10'd 210: cos = 10'd653;
		10'd 211: cos = 10'd650;
		10'd 212: cos = 10'd647;
		10'd 213: cos = 10'd644;
		10'd 214: cos = 10'd641;
		10'd 215: cos = 10'd638;
		10'd 216: cos = 10'd635;
		10'd 217: cos = 10'd632;
		10'd 218: cos = 10'd629;
		10'd 219: cos = 10'd626;
		10'd 220: cos = 10'd623;
		10'd 221: cos = 10'd620;
		10'd 222: cos = 10'd617;
		10'd 223: cos = 10'd614;
		10'd 224: cos = 10'd611;
		10'd 225: cos = 10'd608;
		10'd 226: cos = 10'd605;
		10'd 227: cos = 10'd602;
		10'd 228: cos = 10'd598;
		10'd 229: cos = 10'd595;
		10'd 230: cos = 10'd592;
		10'd 231: cos = 10'd589;
		10'd 232: cos = 10'd586;
		10'd 233: cos = 10'd583;
		10'd 234: cos = 10'd580;
		10'd 235: cos = 10'd577;
		10'd 236: cos = 10'd574;
		10'd 237: cos = 10'd570;
		10'd 238: cos = 10'd567;
		10'd 239: cos = 10'd564;
		10'd 240: cos = 10'd561;
		10'd 241: cos = 10'd558;
		10'd 242: cos = 10'd555;
		10'd 243: cos = 10'd552;
		10'd 244: cos = 10'd549;
		10'd 245: cos = 10'd545;
		10'd 246: cos = 10'd542;
		10'd 247: cos = 10'd539;
		10'd 248: cos = 10'd536;
		10'd 249: cos = 10'd533;
		10'd 250: cos = 10'd530;
		10'd 251: cos = 10'd527;
		10'd 252: cos = 10'd524;
		10'd 253: cos = 10'd520;
		10'd 254: cos = 10'd517;
		10'd 255: cos = 10'd514;
		10'd 256: cos = 10'd511;
		10'd 257: cos = 10'd508;
		10'd 258: cos = 10'd505;
		10'd 259: cos = 10'd502;
		10'd 260: cos = 10'd498;
		10'd 261: cos = 10'd495;
		10'd 262: cos = 10'd492;
		10'd 263: cos = 10'd489;
		10'd 264: cos = 10'd486;
		10'd 265: cos = 10'd483;
		10'd 266: cos = 10'd480;
		10'd 267: cos = 10'd477;
		10'd 268: cos = 10'd473;
		10'd 269: cos = 10'd470;
		10'd 270: cos = 10'd467;
		10'd 271: cos = 10'd464;
		10'd 272: cos = 10'd461;
		10'd 273: cos = 10'd458;
		10'd 274: cos = 10'd455;
		10'd 275: cos = 10'd452;
		10'd 276: cos = 10'd448;
		10'd 277: cos = 10'd445;
		10'd 278: cos = 10'd442;
		10'd 279: cos = 10'd439;
		10'd 280: cos = 10'd436;
		10'd 281: cos = 10'd433;
		10'd 282: cos = 10'd430;
		10'd 283: cos = 10'd427;
		10'd 284: cos = 10'd424;
		10'd 285: cos = 10'd420;
		10'd 286: cos = 10'd417;
		10'd 287: cos = 10'd414;
		10'd 288: cos = 10'd411;
		10'd 289: cos = 10'd408;
		10'd 290: cos = 10'd405;
		10'd 291: cos = 10'd402;
		10'd 292: cos = 10'd399;
		10'd 293: cos = 10'd396;
		10'd 294: cos = 10'd393;
		10'd 295: cos = 10'd390;
		10'd 296: cos = 10'd387;
		10'd 297: cos = 10'd384;
		10'd 298: cos = 10'd381;
		10'd 299: cos = 10'd378;
		10'd 300: cos = 10'd375;
		10'd 301: cos = 10'd372;
		10'd 302: cos = 10'd369;
		10'd 303: cos = 10'd366;
		10'd 304: cos = 10'd363;
		10'd 305: cos = 10'd360;
		10'd 306: cos = 10'd357;
		10'd 307: cos = 10'd354;
		10'd 308: cos = 10'd351;
		10'd 309: cos = 10'd348;
		10'd 310: cos = 10'd345;
		10'd 311: cos = 10'd342;
		10'd 312: cos = 10'd339;
		10'd 313: cos = 10'd336;
		10'd 314: cos = 10'd333;
		10'd 315: cos = 10'd330;
		10'd 316: cos = 10'd327;
		10'd 317: cos = 10'd324;
		10'd 318: cos = 10'd321;
		10'd 319: cos = 10'd318;
		10'd 320: cos = 10'd315;
		10'd 321: cos = 10'd312;
		10'd 322: cos = 10'd309;
		10'd 323: cos = 10'd307;
		10'd 324: cos = 10'd304;
		10'd 325: cos = 10'd301;
		10'd 326: cos = 10'd298;
		10'd 327: cos = 10'd295;
		10'd 328: cos = 10'd292;
		10'd 329: cos = 10'd289;
		10'd 330: cos = 10'd287;
		10'd 331: cos = 10'd284;
		10'd 332: cos = 10'd281;
		10'd 333: cos = 10'd278;
		10'd 334: cos = 10'd275;
		10'd 335: cos = 10'd273;
		10'd 336: cos = 10'd270;
		10'd 337: cos = 10'd267;
		10'd 338: cos = 10'd264;
		10'd 339: cos = 10'd262;
		10'd 340: cos = 10'd259;
		10'd 341: cos = 10'd256;
		10'd 342: cos = 10'd253;
		10'd 343: cos = 10'd251;
		10'd 344: cos = 10'd248;
		10'd 345: cos = 10'd245;
		10'd 346: cos = 10'd243;
		10'd 347: cos = 10'd240;
		10'd 348: cos = 10'd237;
		10'd 349: cos = 10'd235;
		10'd 350: cos = 10'd232;
		10'd 351: cos = 10'd229;
		10'd 352: cos = 10'd227;
		10'd 353: cos = 10'd224;
		10'd 354: cos = 10'd222;
		10'd 355: cos = 10'd219;
		10'd 356: cos = 10'd216;
		10'd 357: cos = 10'd214;
		10'd 358: cos = 10'd211;
		10'd 359: cos = 10'd209;
		10'd 360: cos = 10'd206;
		10'd 361: cos = 10'd204;
		10'd 362: cos = 10'd201;
		10'd 363: cos = 10'd199;
		10'd 364: cos = 10'd196;
		10'd 365: cos = 10'd194;
		10'd 366: cos = 10'd191;
		10'd 367: cos = 10'd189;
		10'd 368: cos = 10'd187;
		10'd 369: cos = 10'd184;
		10'd 370: cos = 10'd182;
		10'd 371: cos = 10'd179;
		10'd 372: cos = 10'd177;
		10'd 373: cos = 10'd175;
		10'd 374: cos = 10'd172;
		10'd 375: cos = 10'd170;
		10'd 376: cos = 10'd167;
		10'd 377: cos = 10'd165;
		10'd 378: cos = 10'd163;
		10'd 379: cos = 10'd161;
		10'd 380: cos = 10'd158;
		10'd 381: cos = 10'd156;
		10'd 382: cos = 10'd154;
		10'd 383: cos = 10'd152;
		10'd 384: cos = 10'd149;
		10'd 385: cos = 10'd147;
		10'd 386: cos = 10'd145;
		10'd 387: cos = 10'd143;
		10'd 388: cos = 10'd141;
		10'd 389: cos = 10'd138;
		10'd 390: cos = 10'd136;
		10'd 391: cos = 10'd134;
		10'd 392: cos = 10'd132;
		10'd 393: cos = 10'd130;
		10'd 394: cos = 10'd128;
		10'd 395: cos = 10'd126;
		10'd 396: cos = 10'd124;
		10'd 397: cos = 10'd122;
		10'd 398: cos = 10'd120;
		10'd 399: cos = 10'd118;
		10'd 400: cos = 10'd116;
		10'd 401: cos = 10'd114;
		10'd 402: cos = 10'd112;
		10'd 403: cos = 10'd110;
		10'd 404: cos = 10'd108;
		10'd 405: cos = 10'd106;
		10'd 406: cos = 10'd104;
		10'd 407: cos = 10'd102;
		10'd 408: cos = 10'd100;
		10'd 409: cos = 10'd98;
		10'd 410: cos = 10'd96;
		10'd 411: cos = 10'd95;
		10'd 412: cos = 10'd93;
		10'd 413: cos = 10'd91;
		10'd 414: cos = 10'd89;
		10'd 415: cos = 10'd87;
		10'd 416: cos = 10'd86;
		10'd 417: cos = 10'd84;
		10'd 418: cos = 10'd82;
		10'd 419: cos = 10'd81;
		10'd 420: cos = 10'd79;
		10'd 421: cos = 10'd77;
		10'd 422: cos = 10'd76;
		10'd 423: cos = 10'd74;
		10'd 424: cos = 10'd72;
		10'd 425: cos = 10'd71;
		10'd 426: cos = 10'd69;
		10'd 427: cos = 10'd68;
		10'd 428: cos = 10'd66;
		10'd 429: cos = 10'd64;
		10'd 430: cos = 10'd63;
		10'd 431: cos = 10'd61;
		10'd 432: cos = 10'd60;
		10'd 433: cos = 10'd58;
		10'd 434: cos = 10'd57;
		10'd 435: cos = 10'd56;
		10'd 436: cos = 10'd54;
		10'd 437: cos = 10'd53;
		10'd 438: cos = 10'd51;
		10'd 439: cos = 10'd50;
		10'd 440: cos = 10'd49;
		10'd 441: cos = 10'd47;
		10'd 442: cos = 10'd46;
		10'd 443: cos = 10'd45;
		10'd 444: cos = 10'd43;
		10'd 445: cos = 10'd42;
		10'd 446: cos = 10'd41;
		10'd 447: cos = 10'd40;
		10'd 448: cos = 10'd38;
		10'd 449: cos = 10'd37;
		10'd 450: cos = 10'd36;
		10'd 451: cos = 10'd35;
		10'd 452: cos = 10'd34;
		10'd 453: cos = 10'd33;
		10'd 454: cos = 10'd32;
		10'd 455: cos = 10'd30;
		10'd 456: cos = 10'd29;
		10'd 457: cos = 10'd28;
		10'd 458: cos = 10'd27;
		10'd 459: cos = 10'd26;
		10'd 460: cos = 10'd25;
		10'd 461: cos = 10'd24;
		10'd 462: cos = 10'd23;
		10'd 463: cos = 10'd22;
		10'd 464: cos = 10'd22;
		10'd 465: cos = 10'd21;
		10'd 466: cos = 10'd20;
		10'd 467: cos = 10'd19;
		10'd 468: cos = 10'd18;
		10'd 469: cos = 10'd17;
		10'd 470: cos = 10'd16;
		10'd 471: cos = 10'd16;
		10'd 472: cos = 10'd15;
		10'd 473: cos = 10'd14;
		10'd 474: cos = 10'd13;
		10'd 475: cos = 10'd13;
		10'd 476: cos = 10'd12;
		10'd 477: cos = 10'd11;
		10'd 478: cos = 10'd11;
		10'd 479: cos = 10'd10;
		10'd 480: cos = 10'd9;
		10'd 481: cos = 10'd9;
		10'd 482: cos = 10'd8;
		10'd 483: cos = 10'd8;
		10'd 484: cos = 10'd7;
		10'd 485: cos = 10'd7;
		10'd 486: cos = 10'd6;
		10'd 487: cos = 10'd6;
		10'd 488: cos = 10'd5;
		10'd 489: cos = 10'd5;
		10'd 490: cos = 10'd4;
		10'd 491: cos = 10'd4;
		10'd 492: cos = 10'd3;
		10'd 493: cos = 10'd3;
		10'd 494: cos = 10'd3;
		10'd 495: cos = 10'd2;
		10'd 496: cos = 10'd2;
		10'd 497: cos = 10'd2;
		10'd 498: cos = 10'd1;
		10'd 499: cos = 10'd1;
		10'd 500: cos = 10'd1;
		10'd 501: cos = 10'd1;
		10'd 502: cos = 10'd0;
		10'd 503: cos = 10'd0;
		10'd 504: cos = 10'd0;
		10'd 505: cos = 10'd0;
		10'd 506: cos = 10'd0;
		10'd 507: cos = 10'd0;
		10'd 508: cos = 10'd0;
		10'd 509: cos = 10'd0;
		10'd 510: cos = 10'd0;
		10'd 511: cos = 10'd0;
		10'd 512: cos = 10'd0;
		10'd 513: cos = 10'd0;
		10'd 514: cos = 10'd0;
		10'd 515: cos = 10'd0;
		10'd 516: cos = 10'd0;
		10'd 517: cos = 10'd0;
		10'd 518: cos = 10'd0;
		10'd 519: cos = 10'd0;
		10'd 520: cos = 10'd0;
		10'd 521: cos = 10'd0;
		10'd 522: cos = 10'd0;
		10'd 523: cos = 10'd1;
		10'd 524: cos = 10'd1;
		10'd 525: cos = 10'd1;
		10'd 526: cos = 10'd1;
		10'd 527: cos = 10'd2;
		10'd 528: cos = 10'd2;
		10'd 529: cos = 10'd2;
		10'd 530: cos = 10'd3;
		10'd 531: cos = 10'd3;
		10'd 532: cos = 10'd3;
		10'd 533: cos = 10'd4;
		10'd 534: cos = 10'd4;
		10'd 535: cos = 10'd5;
		10'd 536: cos = 10'd5;
		10'd 537: cos = 10'd6;
		10'd 538: cos = 10'd6;
		10'd 539: cos = 10'd7;
		10'd 540: cos = 10'd7;
		10'd 541: cos = 10'd8;
		10'd 542: cos = 10'd8;
		10'd 543: cos = 10'd9;
		10'd 544: cos = 10'd9;
		10'd 545: cos = 10'd10;
		10'd 546: cos = 10'd11;
		10'd 547: cos = 10'd11;
		10'd 548: cos = 10'd12;
		10'd 549: cos = 10'd13;
		10'd 550: cos = 10'd13;
		10'd 551: cos = 10'd14;
		10'd 552: cos = 10'd15;
		10'd 553: cos = 10'd16;
		10'd 554: cos = 10'd16;
		10'd 555: cos = 10'd17;
		10'd 556: cos = 10'd18;
		10'd 557: cos = 10'd19;
		10'd 558: cos = 10'd20;
		10'd 559: cos = 10'd21;
		10'd 560: cos = 10'd22;
		10'd 561: cos = 10'd22;
		10'd 562: cos = 10'd23;
		10'd 563: cos = 10'd24;
		10'd 564: cos = 10'd25;
		10'd 565: cos = 10'd26;
		10'd 566: cos = 10'd27;
		10'd 567: cos = 10'd28;
		10'd 568: cos = 10'd29;
		10'd 569: cos = 10'd30;
		10'd 570: cos = 10'd32;
		10'd 571: cos = 10'd33;
		10'd 572: cos = 10'd34;
		10'd 573: cos = 10'd35;
		10'd 574: cos = 10'd36;
		10'd 575: cos = 10'd37;
		10'd 576: cos = 10'd38;
		10'd 577: cos = 10'd40;
		10'd 578: cos = 10'd41;
		10'd 579: cos = 10'd42;
		10'd 580: cos = 10'd43;
		10'd 581: cos = 10'd45;
		10'd 582: cos = 10'd46;
		10'd 583: cos = 10'd47;
		10'd 584: cos = 10'd49;
		10'd 585: cos = 10'd50;
		10'd 586: cos = 10'd51;
		10'd 587: cos = 10'd53;
		10'd 588: cos = 10'd54;
		10'd 589: cos = 10'd56;
		10'd 590: cos = 10'd57;
		10'd 591: cos = 10'd58;
		10'd 592: cos = 10'd60;
		10'd 593: cos = 10'd61;
		10'd 594: cos = 10'd63;
		10'd 595: cos = 10'd64;
		10'd 596: cos = 10'd66;
		10'd 597: cos = 10'd68;
		10'd 598: cos = 10'd69;
		10'd 599: cos = 10'd71;
		10'd 600: cos = 10'd72;
		10'd 601: cos = 10'd74;
		10'd 602: cos = 10'd76;
		10'd 603: cos = 10'd77;
		10'd 604: cos = 10'd79;
		10'd 605: cos = 10'd81;
		10'd 606: cos = 10'd82;
		10'd 607: cos = 10'd84;
		10'd 608: cos = 10'd86;
		10'd 609: cos = 10'd87;
		10'd 610: cos = 10'd89;
		10'd 611: cos = 10'd91;
		10'd 612: cos = 10'd93;
		10'd 613: cos = 10'd95;
		10'd 614: cos = 10'd96;
		10'd 615: cos = 10'd98;
		10'd 616: cos = 10'd100;
		10'd 617: cos = 10'd102;
		10'd 618: cos = 10'd104;
		10'd 619: cos = 10'd106;
		10'd 620: cos = 10'd108;
		10'd 621: cos = 10'd110;
		10'd 622: cos = 10'd112;
		10'd 623: cos = 10'd114;
		10'd 624: cos = 10'd116;
		10'd 625: cos = 10'd118;
		10'd 626: cos = 10'd120;
		10'd 627: cos = 10'd122;
		10'd 628: cos = 10'd124;
		10'd 629: cos = 10'd126;
		10'd 630: cos = 10'd128;
		10'd 631: cos = 10'd130;
		10'd 632: cos = 10'd132;
		10'd 633: cos = 10'd134;
		10'd 634: cos = 10'd136;
		10'd 635: cos = 10'd138;
		10'd 636: cos = 10'd141;
		10'd 637: cos = 10'd143;
		10'd 638: cos = 10'd145;
		10'd 639: cos = 10'd147;
		10'd 640: cos = 10'd149;
		10'd 641: cos = 10'd152;
		10'd 642: cos = 10'd154;
		10'd 643: cos = 10'd156;
		10'd 644: cos = 10'd158;
		10'd 645: cos = 10'd161;
		10'd 646: cos = 10'd163;
		10'd 647: cos = 10'd165;
		10'd 648: cos = 10'd167;
		10'd 649: cos = 10'd170;
		10'd 650: cos = 10'd172;
		10'd 651: cos = 10'd175;
		10'd 652: cos = 10'd177;
		10'd 653: cos = 10'd179;
		10'd 654: cos = 10'd182;
		10'd 655: cos = 10'd184;
		10'd 656: cos = 10'd187;
		10'd 657: cos = 10'd189;
		10'd 658: cos = 10'd191;
		10'd 659: cos = 10'd194;
		10'd 660: cos = 10'd196;
		10'd 661: cos = 10'd199;
		10'd 662: cos = 10'd201;
		10'd 663: cos = 10'd204;
		10'd 664: cos = 10'd206;
		10'd 665: cos = 10'd209;
		10'd 666: cos = 10'd211;
		10'd 667: cos = 10'd214;
		10'd 668: cos = 10'd216;
		10'd 669: cos = 10'd219;
		10'd 670: cos = 10'd222;
		10'd 671: cos = 10'd224;
		10'd 672: cos = 10'd227;
		10'd 673: cos = 10'd229;
		10'd 674: cos = 10'd232;
		10'd 675: cos = 10'd235;
		10'd 676: cos = 10'd237;
		10'd 677: cos = 10'd240;
		10'd 678: cos = 10'd243;
		10'd 679: cos = 10'd245;
		10'd 680: cos = 10'd248;
		10'd 681: cos = 10'd251;
		10'd 682: cos = 10'd253;
		10'd 683: cos = 10'd256;
		10'd 684: cos = 10'd259;
		10'd 685: cos = 10'd262;
		10'd 686: cos = 10'd264;
		10'd 687: cos = 10'd267;
		10'd 688: cos = 10'd270;
		10'd 689: cos = 10'd273;
		10'd 690: cos = 10'd275;
		10'd 691: cos = 10'd278;
		10'd 692: cos = 10'd281;
		10'd 693: cos = 10'd284;
		10'd 694: cos = 10'd287;
		10'd 695: cos = 10'd289;
		10'd 696: cos = 10'd292;
		10'd 697: cos = 10'd295;
		10'd 698: cos = 10'd298;
		10'd 699: cos = 10'd301;
		10'd 700: cos = 10'd304;
		10'd 701: cos = 10'd307;
		10'd 702: cos = 10'd309;
		10'd 703: cos = 10'd312;
		10'd 704: cos = 10'd315;
		10'd 705: cos = 10'd318;
		10'd 706: cos = 10'd321;
		10'd 707: cos = 10'd324;
		10'd 708: cos = 10'd327;
		10'd 709: cos = 10'd330;
		10'd 710: cos = 10'd333;
		10'd 711: cos = 10'd336;
		10'd 712: cos = 10'd339;
		10'd 713: cos = 10'd342;
		10'd 714: cos = 10'd345;
		10'd 715: cos = 10'd348;
		10'd 716: cos = 10'd351;
		10'd 717: cos = 10'd354;
		10'd 718: cos = 10'd357;
		10'd 719: cos = 10'd360;
		10'd 720: cos = 10'd363;
		10'd 721: cos = 10'd366;
		10'd 722: cos = 10'd369;
		10'd 723: cos = 10'd372;
		10'd 724: cos = 10'd375;
		10'd 725: cos = 10'd378;
		10'd 726: cos = 10'd381;
		10'd 727: cos = 10'd384;
		10'd 728: cos = 10'd387;
		10'd 729: cos = 10'd390;
		10'd 730: cos = 10'd393;
		10'd 731: cos = 10'd396;
		10'd 732: cos = 10'd399;
		10'd 733: cos = 10'd402;
		10'd 734: cos = 10'd405;
		10'd 735: cos = 10'd408;
		10'd 736: cos = 10'd411;
		10'd 737: cos = 10'd414;
		10'd 738: cos = 10'd417;
		10'd 739: cos = 10'd420;
		10'd 740: cos = 10'd424;
		10'd 741: cos = 10'd427;
		10'd 742: cos = 10'd430;
		10'd 743: cos = 10'd433;
		10'd 744: cos = 10'd436;
		10'd 745: cos = 10'd439;
		10'd 746: cos = 10'd442;
		10'd 747: cos = 10'd445;
		10'd 748: cos = 10'd448;
		10'd 749: cos = 10'd452;
		10'd 750: cos = 10'd455;
		10'd 751: cos = 10'd458;
		10'd 752: cos = 10'd461;
		10'd 753: cos = 10'd464;
		10'd 754: cos = 10'd467;
		10'd 755: cos = 10'd470;
		10'd 756: cos = 10'd473;
		10'd 757: cos = 10'd477;
		10'd 758: cos = 10'd480;
		10'd 759: cos = 10'd483;
		10'd 760: cos = 10'd486;
		10'd 761: cos = 10'd489;
		10'd 762: cos = 10'd492;
		10'd 763: cos = 10'd495;
		10'd 764: cos = 10'd498;
		10'd 765: cos = 10'd502;
		10'd 766: cos = 10'd505;
		10'd 767: cos = 10'd508;
		10'd 768: cos = 10'd511;
		10'd 769: cos = 10'd514;
		10'd 770: cos = 10'd517;
		10'd 771: cos = 10'd520;
		10'd 772: cos = 10'd524;
		10'd 773: cos = 10'd527;
		10'd 774: cos = 10'd530;
		10'd 775: cos = 10'd533;
		10'd 776: cos = 10'd536;
		10'd 777: cos = 10'd539;
		10'd 778: cos = 10'd542;
		10'd 779: cos = 10'd545;
		10'd 780: cos = 10'd549;
		10'd 781: cos = 10'd552;
		10'd 782: cos = 10'd555;
		10'd 783: cos = 10'd558;
		10'd 784: cos = 10'd561;
		10'd 785: cos = 10'd564;
		10'd 786: cos = 10'd567;
		10'd 787: cos = 10'd570;
		10'd 788: cos = 10'd574;
		10'd 789: cos = 10'd577;
		10'd 790: cos = 10'd580;
		10'd 791: cos = 10'd583;
		10'd 792: cos = 10'd586;
		10'd 793: cos = 10'd589;
		10'd 794: cos = 10'd592;
		10'd 795: cos = 10'd595;
		10'd 796: cos = 10'd598;
		10'd 797: cos = 10'd602;
		10'd 798: cos = 10'd605;
		10'd 799: cos = 10'd608;
		10'd 800: cos = 10'd611;
		10'd 801: cos = 10'd614;
		10'd 802: cos = 10'd617;
		10'd 803: cos = 10'd620;
		10'd 804: cos = 10'd623;
		10'd 805: cos = 10'd626;
		10'd 806: cos = 10'd629;
		10'd 807: cos = 10'd632;
		10'd 808: cos = 10'd635;
		10'd 809: cos = 10'd638;
		10'd 810: cos = 10'd641;
		10'd 811: cos = 10'd644;
		10'd 812: cos = 10'd647;
		10'd 813: cos = 10'd650;
		10'd 814: cos = 10'd653;
		10'd 815: cos = 10'd656;
		10'd 816: cos = 10'd659;
		10'd 817: cos = 10'd662;
		10'd 818: cos = 10'd665;
		10'd 819: cos = 10'd668;
		10'd 820: cos = 10'd671;
		10'd 821: cos = 10'd674;
		10'd 822: cos = 10'd677;
		10'd 823: cos = 10'd680;
		10'd 824: cos = 10'd683;
		10'd 825: cos = 10'd686;
		10'd 826: cos = 10'd689;
		10'd 827: cos = 10'd692;
		10'd 828: cos = 10'd695;
		10'd 829: cos = 10'd698;
		10'd 830: cos = 10'd701;
		10'd 831: cos = 10'd704;
		10'd 832: cos = 10'd707;
		10'd 833: cos = 10'd710;
		10'd 834: cos = 10'd713;
		10'd 835: cos = 10'd715;
		10'd 836: cos = 10'd718;
		10'd 837: cos = 10'd721;
		10'd 838: cos = 10'd724;
		10'd 839: cos = 10'd727;
		10'd 840: cos = 10'd730;
		10'd 841: cos = 10'd733;
		10'd 842: cos = 10'd735;
		10'd 843: cos = 10'd738;
		10'd 844: cos = 10'd741;
		10'd 845: cos = 10'd744;
		10'd 846: cos = 10'd747;
		10'd 847: cos = 10'd749;
		10'd 848: cos = 10'd752;
		10'd 849: cos = 10'd755;
		10'd 850: cos = 10'd758;
		10'd 851: cos = 10'd760;
		10'd 852: cos = 10'd763;
		10'd 853: cos = 10'd766;
		10'd 854: cos = 10'd769;
		10'd 855: cos = 10'd771;
		10'd 856: cos = 10'd774;
		10'd 857: cos = 10'd777;
		10'd 858: cos = 10'd779;
		10'd 859: cos = 10'd782;
		10'd 860: cos = 10'd785;
		10'd 861: cos = 10'd787;
		10'd 862: cos = 10'd790;
		10'd 863: cos = 10'd793;
		10'd 864: cos = 10'd795;
		10'd 865: cos = 10'd798;
		10'd 866: cos = 10'd800;
		10'd 867: cos = 10'd803;
		10'd 868: cos = 10'd806;
		10'd 869: cos = 10'd808;
		10'd 870: cos = 10'd811;
		10'd 871: cos = 10'd813;
		10'd 872: cos = 10'd816;
		10'd 873: cos = 10'd818;
		10'd 874: cos = 10'd821;
		10'd 875: cos = 10'd823;
		10'd 876: cos = 10'd826;
		10'd 877: cos = 10'd828;
		10'd 878: cos = 10'd831;
		10'd 879: cos = 10'd833;
		10'd 880: cos = 10'd835;
		10'd 881: cos = 10'd838;
		10'd 882: cos = 10'd840;
		10'd 883: cos = 10'd843;
		10'd 884: cos = 10'd845;
		10'd 885: cos = 10'd847;
		10'd 886: cos = 10'd850;
		10'd 887: cos = 10'd852;
		10'd 888: cos = 10'd855;
		10'd 889: cos = 10'd857;
		10'd 890: cos = 10'd859;
		10'd 891: cos = 10'd861;
		10'd 892: cos = 10'd864;
		10'd 893: cos = 10'd866;
		10'd 894: cos = 10'd868;
		10'd 895: cos = 10'd870;
		10'd 896: cos = 10'd873;
		10'd 897: cos = 10'd875;
		10'd 898: cos = 10'd877;
		10'd 899: cos = 10'd879;
		10'd 900: cos = 10'd881;
		10'd 901: cos = 10'd884;
		10'd 902: cos = 10'd886;
		10'd 903: cos = 10'd888;
		10'd 904: cos = 10'd890;
		10'd 905: cos = 10'd892;
		10'd 906: cos = 10'd894;
		10'd 907: cos = 10'd896;
		10'd 908: cos = 10'd898;
		10'd 909: cos = 10'd900;
		10'd 910: cos = 10'd902;
		10'd 911: cos = 10'd904;
		10'd 912: cos = 10'd906;
		10'd 913: cos = 10'd908;
		10'd 914: cos = 10'd910;
		10'd 915: cos = 10'd912;
		10'd 916: cos = 10'd914;
		10'd 917: cos = 10'd916;
		10'd 918: cos = 10'd918;
		10'd 919: cos = 10'd920;
		10'd 920: cos = 10'd922;
		10'd 921: cos = 10'd924;
		10'd 922: cos = 10'd926;
		10'd 923: cos = 10'd927;
		10'd 924: cos = 10'd929;
		10'd 925: cos = 10'd931;
		10'd 926: cos = 10'd933;
		10'd 927: cos = 10'd935;
		10'd 928: cos = 10'd936;
		10'd 929: cos = 10'd938;
		10'd 930: cos = 10'd940;
		10'd 931: cos = 10'd941;
		10'd 932: cos = 10'd943;
		10'd 933: cos = 10'd945;
		10'd 934: cos = 10'd946;
		10'd 935: cos = 10'd948;
		10'd 936: cos = 10'd950;
		10'd 937: cos = 10'd951;
		10'd 938: cos = 10'd953;
		10'd 939: cos = 10'd954;
		10'd 940: cos = 10'd956;
		10'd 941: cos = 10'd958;
		10'd 942: cos = 10'd959;
		10'd 943: cos = 10'd961;
		10'd 944: cos = 10'd962;
		10'd 945: cos = 10'd964;
		10'd 946: cos = 10'd965;
		10'd 947: cos = 10'd966;
		10'd 948: cos = 10'd968;
		10'd 949: cos = 10'd969;
		10'd 950: cos = 10'd971;
		10'd 951: cos = 10'd972;
		10'd 952: cos = 10'd973;
		10'd 953: cos = 10'd975;
		10'd 954: cos = 10'd976;
		10'd 955: cos = 10'd977;
		10'd 956: cos = 10'd979;
		10'd 957: cos = 10'd980;
		10'd 958: cos = 10'd981;
		10'd 959: cos = 10'd982;
		10'd 960: cos = 10'd984;
		10'd 961: cos = 10'd985;
		10'd 962: cos = 10'd986;
		10'd 963: cos = 10'd987;
		10'd 964: cos = 10'd988;
		10'd 965: cos = 10'd989;
		10'd 966: cos = 10'd990;
		10'd 967: cos = 10'd992;
		10'd 968: cos = 10'd993;
		10'd 969: cos = 10'd994;
		10'd 970: cos = 10'd995;
		10'd 971: cos = 10'd996;
		10'd 972: cos = 10'd997;
		10'd 973: cos = 10'd998;
		10'd 974: cos = 10'd999;
		10'd 975: cos = 10'd1000;
		10'd 976: cos = 10'd1000;
		10'd 977: cos = 10'd1001;
		10'd 978: cos = 10'd1002;
		10'd 979: cos = 10'd1003;
		10'd 980: cos = 10'd1004;
		10'd 981: cos = 10'd1005;
		10'd 982: cos = 10'd1006;
		10'd 983: cos = 10'd1006;
		10'd 984: cos = 10'd1007;
		10'd 985: cos = 10'd1008;
		10'd 986: cos = 10'd1009;
		10'd 987: cos = 10'd1009;
		10'd 988: cos = 10'd1010;
		10'd 989: cos = 10'd1011;
		10'd 990: cos = 10'd1011;
		10'd 991: cos = 10'd1012;
		10'd 992: cos = 10'd1013;
		10'd 993: cos = 10'd1013;
		10'd 994: cos = 10'd1014;
		10'd 995: cos = 10'd1014;
		10'd 996: cos = 10'd1015;
		10'd 997: cos = 10'd1015;
		10'd 998: cos = 10'd1016;
		10'd 999: cos = 10'd1016;
		10'd1000: cos = 10'd1017;
		10'd1001: cos = 10'd1017;
		10'd1002: cos = 10'd1018;
		10'd1003: cos = 10'd1018;
		10'd1004: cos = 10'd1019;
		10'd1005: cos = 10'd1019;
		10'd1006: cos = 10'd1019;
		10'd1007: cos = 10'd1020;
		10'd1008: cos = 10'd1020;
		10'd1009: cos = 10'd1020;
		10'd1010: cos = 10'd1021;
		10'd1011: cos = 10'd1021;
		10'd1012: cos = 10'd1021;
		10'd1013: cos = 10'd1021;
		10'd1014: cos = 10'd1022;
		10'd1015: cos = 10'd1022;
		10'd1016: cos = 10'd1022;
		10'd1017: cos = 10'd1022;
		10'd1018: cos = 10'd1022;
		10'd1019: cos = 10'd1022;
		10'd1020: cos = 10'd1022;
		10'd1021: cos = 10'd1022;
		10'd1022: cos = 10'd1022;
		default:  cos = 10'd1022;
		endcase
	end
endfunction

endmodule
