module i2c_slave (
	input	wire sda,
	input	wire scl,
	output wire [7:0] led
);

